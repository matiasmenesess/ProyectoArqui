module datapath (
);

endmodule
