module datapath (
	
);

	
endmodule
